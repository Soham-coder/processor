//Global defines goes here

`define WORD_SIZE 32
`define NUMBER_OF_REGISTERS 32
`define OPERATION_TYPE_WIDTH 2

`define NUMBER_OF_PC_REGISTERS 256
`define OPCODE_WIDTH 5